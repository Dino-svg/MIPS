module SUM( 
    input data,
    output DataOut
);

    assign DataOut= 4 + data;
	
endmodule
