module SUM( 
    input data,
    output dataOut
);

    dataOut= 4 + data;
	
endmodule
